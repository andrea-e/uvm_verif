`ifndef RESET_SEQ_LIB_SV
 `define RESET_SEQ_LIB_SV

 `include "sequences/reset_base_seq.sv"
 `include "sequences/reset_seq.sv"

`endif
