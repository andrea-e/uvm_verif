`ifndef APB_SLAVE_SEQ_LIB_SV
 `define APB_SLAVE_SEQ_LIB_SV

 `include "slave/sequences/apb_slave_base_seq.sv"
 `include "slave/sequences/apb_slave_simple_seq.sv"

`endif
