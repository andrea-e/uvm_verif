`ifndef I2C_SLAVE_SEQ_LIB_SV
 `define I2C_SLAVE_SEQ_LIB_SV

 `include "slave/sequences/i2c_slave_base_seq.sv"
 `include "slave/sequences/i2c_slave_simple_seq.sv"

`endif
