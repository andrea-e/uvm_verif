`ifndef RESET_IF_SV
 `define RESET_IF_SV

interface reset_if (input clk, output logic reset);

endinterface : reset_if

`endif
