`ifndef I2C_MASTER_SEQ_LIB_SV
 `define I2C_MASTER_SEQ_LIB_SV

 `include "master/sequences/i2c_master_base_seq.sv"
 `include "master/sequences/i2c_master_simple_seq.sv"

`endif
