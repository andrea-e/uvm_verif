`ifndef APB_TYPES_SV
 `define APB_TYPES_SV

typedef enum {
              APB_READ = 0,
              APB_WRITE = 1
              } apb_direction_enum;

`endif
