`ifndef I2C_TEST_LIB_SV
 `define I2C_TEST_LIB_SV

 `include "i2c_test_base.sv"
 `include "i2c_test_simple.sv"

`endif
