`ifndef RESET_PKG_SV
 `define RESET_PKG_SV

package reset_pkg;

   import uvm_pkg::*;
 `include "uvm_macros.svh"

 `include "reset_config.sv"
 `include "reset_seq_item.sv"
 `include "reset_driver.sv"
 `include "reset_monitor.sv"
 `include "reset_agent.sv"
 `include "sequences/reset_seq_lib.sv"

endpackage : reset_pkg

 `include "reset_if.sv"

`endif
