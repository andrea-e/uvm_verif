`ifndef CALC_SEQ_LIB_SV
 `define CALC_SEQ_LIB_SV

 `include "sequences/v8_calc_base_seq.sv"
 `include "sequences/v8_calc_simple_seq.sv"

`endif
