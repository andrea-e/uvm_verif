`ifndef APB_MASTER_SEQ_LIB_SV
 `define APB_MASTER_SEQ_LIB_SV

 `include "master/sequences/apb_master_base_seq.sv"
 `include "master/sequences/apb_master_simple_seq.sv"
 `include "master/sequences/apb_master_read_seq.sv"
 `include "master/sequences/apb_master_write_seq.sv"
 `include "master/sequences/apb_master_read_all_seq.sv"
 `include "master/sequences/apb_master_write_all_seq.sv"
 `include "master/sequences/apb_master_read_after_write_seq.sv"

`endif
