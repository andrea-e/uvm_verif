`ifndef TEST_LIB_SV
 `define TEST_LIB_SV

 `include "tests/v10_test_base.sv"
 `include "tests/v10_test_simple.sv"
 `include "tests/v10_test_simple_2.sv"

`endif
