`ifndef APB_TEST_LIB_SV
 `define APB_TEST_LIB_SV

 `include "apb_test_base.sv"
 `include "apb_test_simple.sv"

`endif
