class calc_config extends uvm_object;

   uvm_active_passive_enum is_active = UVM_ACTIVE;

   `uvm_object_utils_begin (calc_config)
      `uvm_field_enum(uvm_active_passive_enum, is_active, UVM_DEFAULT)
   `uvm_object_utils_end

   function new(string name = "calc_config");
      super.new(name);
   endfunction

endclass : calc_config
