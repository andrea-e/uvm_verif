`ifndef MEMORY_PKG_SV
 `define MEMORY_PKG_SV

package memory_pkg;

 `include "v2_tr.sv"
 `include "v2_driver.sv"

endpackage : memory_pkg

`endif
